module mux_4x1_32(output[31:0] o,input[31:0] x0,input[31:0] x1,input[31:0]x2,input[31:0] x3,input s1,input s0);

mux_4x1 m0(o[0],x0[0],x1[0],x2[0],x3[0],s1,s0);
mux_4x1 m1(o[1],x0[1],x1[1],x2[1],x3[1],s1,s0);
mux_4x1 m2(o[2],x0[2],x1[2],x2[2],x3[2],s1,s0);
mux_4x1 m3(o[3],x0[3],x1[3],x2[3],x3[3],s1,s0);
mux_4x1 m4(o[4],x0[4],x1[4],x2[4],x3[4],s1,s0);
mux_4x1 m5(o[5],x0[5],x1[5],x2[5],x3[5],s1,s0);
mux_4x1 m6(o[6],x0[6],x1[6],x2[6],x3[6],s1,s0);
mux_4x1 m7(o[7],x0[7],x1[7],x2[7],x3[7],s1,s0);
mux_4x1 m8(o[8],x0[8],x1[8],x2[8],x3[8],s1,s0);
mux_4x1 m9(o[9],x0[9],x1[9],x2[9],x3[9],s1,s0);
mux_4x1 m10(o[10],x0[10],x1[10],x2[10],x3[10],s1,s0);
mux_4x1 m11(o[11],x0[11],x1[11],x2[11],x3[11],s1,s0);
mux_4x1 m12(o[12],x0[12],x1[12],x2[12],x3[12],s1,s0);
mux_4x1 m13(o[13],x0[13],x1[13],x2[13],x3[13],s1,s0);
mux_4x1 m14(o[14],x0[14],x1[14],x2[14],x3[14],s1,s0);
mux_4x1 m15(o[15],x0[15],x1[15],x2[15],x3[15],s1,s0);
mux_4x1 m16(o[16],x0[16],x1[16],x2[16],x3[16],s1,s0);
mux_4x1 m17(o[17],x0[17],x1[17],x2[17],x3[17],s1,s0);
mux_4x1 m18(o[18],x0[18],x1[18],x2[18],x3[18],s1,s0);
mux_4x1 m19(o[19],x0[19],x1[19],x2[19],x3[19],s1,s0);
mux_4x1 m20(o[20],x0[20],x1[20],x2[20],x3[20],s1,s0);
mux_4x1 m21(o[21],x0[21],x1[21],x2[21],x3[21],s1,s0);
mux_4x1 m22(o[22],x0[22],x1[22],x2[22],x3[22],s1,s0);
mux_4x1 m23(o[23],x0[23],x1[23],x2[23],x3[23],s1,s0);
mux_4x1 m24(o[24],x0[24],x1[24],x2[24],x3[24],s1,s0);
mux_4x1 m25(o[25],x0[25],x1[25],x2[25],x3[25],s1,s0);
mux_4x1 m26(o[26],x0[26],x1[26],x2[26],x3[26],s1,s0);
mux_4x1 m27(o[27],x0[27],x1[27],x2[27],x3[27],s1,s0);
mux_4x1 m28(o[28],x0[28],x1[28],x2[28],x3[28],s1,s0);
mux_4x1 m29(o[29],x0[29],x1[29],x2[29],x3[29],s1,s0);
mux_4x1 m30(o[30],x0[30],x1[30],x2[30],x3[30],s1,s0);
mux_4x1 m31(o[31],x0[31],x1[31],x2[31],x3[31],s1,s0);

endmodule