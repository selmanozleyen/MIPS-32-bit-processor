`define DELAY 20
module alu_testbench(); 
reg a, b, carry_in ,op0,op1,op2,lessi;
wire res, carry_out;

alu_1 fatb(res, carry_out, carry_in, a, b ,op2,op1,op0,lessi);

initial begin
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b0;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b0; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b0; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b0 ;op2 = 1'b0;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b0;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b0;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;
lessi=1'b1;a = 1'b1; b = 1'b1; carry_in = 1'b1 ;op2 = 1'b1;op1 = 1'b1;op0 = 1'b1;
#`DELAY;


end
 
initial
begin
$monitor("time = %2d, a =%1b, b=%1b, carry_in=%1b, res=%1b, carry_out=%1b , lessi = %1b opcode =%1b%1b%1b", $time, a, b, carry_in, res, carry_out,lessi,
op2,op1,op0);
end
 
endmodule