module shifter(output[31:0] out,input[31:0] in,input rev,input arithmetic,input[4:0] amt);

wire[31:0] new_in;
mux_2x1 r0(new_in[0],in[0],in[31],rev);
mux_2x1 r1(new_in[1],in[1],in[30],rev);
mux_2x1 r2(new_in[2],in[2],in[29],rev);
mux_2x1 r3(new_in[3],in[3],in[28],rev);
mux_2x1 r4(new_in[4],in[4],in[27],rev);
mux_2x1 r5(new_in[5],in[5],in[26],rev);
mux_2x1 r6(new_in[6],in[6],in[25],rev);
mux_2x1 r7(new_in[7],in[7],in[24],rev);
mux_2x1 r8(new_in[8],in[8],in[23],rev);
mux_2x1 r9(new_in[9],in[9],in[22],rev);
mux_2x1 r10(new_in[10],in[10],in[21],rev);
mux_2x1 r11(new_in[11],in[11],in[20],rev);
mux_2x1 r12(new_in[12],in[12],in[19],rev);
mux_2x1 r13(new_in[13],in[13],in[18],rev);
mux_2x1 r14(new_in[14],in[14],in[17],rev);
mux_2x1 r15(new_in[15],in[15],in[16],rev);
mux_2x1 r16(new_in[16],in[16],in[15],rev);
mux_2x1 r17(new_in[17],in[17],in[14],rev);
mux_2x1 r18(new_in[18],in[18],in[13],rev);
mux_2x1 r19(new_in[19],in[19],in[12],rev);
mux_2x1 r20(new_in[20],in[20],in[11],rev);
mux_2x1 r21(new_in[21],in[21],in[10],rev);
mux_2x1 r22(new_in[22],in[22],in[9],rev);
mux_2x1 r23(new_in[23],in[23],in[8],rev);
mux_2x1 r24(new_in[24],in[24],in[7],rev);
mux_2x1 r25(new_in[25],in[25],in[6],rev);
mux_2x1 r26(new_in[26],in[26],in[5],rev);
mux_2x1 r27(new_in[27],in[27],in[4],rev);
mux_2x1 r28(new_in[28],in[28],in[3],rev);
mux_2x1 r29(new_in[29],in[29],in[2],rev);
mux_2x1 r30(new_in[30],in[30],in[1],rev);
mux_2x1 r31(new_in[31],in[31],in[0],rev);

wire empty;
and a1(empty,arithmetic,new_in[31]);

wire[31:0] layer1,layer2,layer3,layer4,layer5;

mux_2x1 L1_0(layer1[0],new_in[0],new_in[1],amt[0]);
mux_2x1 L1_1(layer1[1],new_in[1],new_in[2],amt[0]);
mux_2x1 L1_2(layer1[2],new_in[2],new_in[3],amt[0]);
mux_2x1 L1_3(layer1[3],new_in[3],new_in[4],amt[0]);
mux_2x1 L1_4(layer1[4],new_in[4],new_in[5],amt[0]);
mux_2x1 L1_5(layer1[5],new_in[5],new_in[6],amt[0]);
mux_2x1 L1_6(layer1[6],new_in[6],new_in[7],amt[0]);
mux_2x1 L1_7(layer1[7],new_in[7],new_in[8],amt[0]);
mux_2x1 L1_8(layer1[8],new_in[8],new_in[9],amt[0]);
mux_2x1 L1_9(layer1[9],new_in[9],new_in[10],amt[0]);
mux_2x1 L1_10(layer1[10],new_in[10],new_in[11],amt[0]);
mux_2x1 L1_11(layer1[11],new_in[11],new_in[12],amt[0]);
mux_2x1 L1_12(layer1[12],new_in[12],new_in[13],amt[0]);
mux_2x1 L1_13(layer1[13],new_in[13],new_in[14],amt[0]);
mux_2x1 L1_14(layer1[14],new_in[14],new_in[15],amt[0]);
mux_2x1 L1_15(layer1[15],new_in[15],new_in[16],amt[0]);
mux_2x1 L1_16(layer1[16],new_in[16],new_in[17],amt[0]);
mux_2x1 L1_17(layer1[17],new_in[17],new_in[18],amt[0]);
mux_2x1 L1_18(layer1[18],new_in[18],new_in[19],amt[0]);
mux_2x1 L1_19(layer1[19],new_in[19],new_in[20],amt[0]);
mux_2x1 L1_20(layer1[20],new_in[20],new_in[21],amt[0]);
mux_2x1 L1_21(layer1[21],new_in[21],new_in[22],amt[0]);
mux_2x1 L1_22(layer1[22],new_in[22],new_in[23],amt[0]);
mux_2x1 L1_23(layer1[23],new_in[23],new_in[24],amt[0]);
mux_2x1 L1_24(layer1[24],new_in[24],new_in[25],amt[0]);
mux_2x1 L1_25(layer1[25],new_in[25],new_in[26],amt[0]);
mux_2x1 L1_26(layer1[26],new_in[26],new_in[27],amt[0]);
mux_2x1 L1_27(layer1[27],new_in[27],new_in[28],amt[0]);
mux_2x1 L1_28(layer1[28],new_in[28],new_in[29],amt[0]);
mux_2x1 L1_29(layer1[29],new_in[29],new_in[30],amt[0]);
mux_2x1 L1_30(layer1[30],new_in[30],new_in[31],amt[0]);
mux_2x1 L1_31(layer1[31],new_in[31],empty,amt[0]);

mux_2x1 L2_0(layer2[0],layer1[0],layer1[2],amt[1]);
mux_2x1 L2_1(layer2[1],layer1[1],layer1[3],amt[1]);
mux_2x1 L2_2(layer2[2],layer1[2],layer1[4],amt[1]);
mux_2x1 L2_3(layer2[3],layer1[3],layer1[5],amt[1]);
mux_2x1 L2_4(layer2[4],layer1[4],layer1[6],amt[1]);
mux_2x1 L2_5(layer2[5],layer1[5],layer1[7],amt[1]);
mux_2x1 L2_6(layer2[6],layer1[6],layer1[8],amt[1]);
mux_2x1 L2_7(layer2[7],layer1[7],layer1[9],amt[1]);
mux_2x1 L2_8(layer2[8],layer1[8],layer1[10],amt[1]);
mux_2x1 L2_9(layer2[9],layer1[9],layer1[11],amt[1]);
mux_2x1 L2_10(layer2[10],layer1[10],layer1[12],amt[1]);
mux_2x1 L2_11(layer2[11],layer1[11],layer1[13],amt[1]);
mux_2x1 L2_12(layer2[12],layer1[12],layer1[14],amt[1]);
mux_2x1 L2_13(layer2[13],layer1[13],layer1[15],amt[1]);
mux_2x1 L2_14(layer2[14],layer1[14],layer1[16],amt[1]);
mux_2x1 L2_15(layer2[15],layer1[15],layer1[17],amt[1]);
mux_2x1 L2_16(layer2[16],layer1[16],layer1[18],amt[1]);
mux_2x1 L2_17(layer2[17],layer1[17],layer1[19],amt[1]);
mux_2x1 L2_18(layer2[18],layer1[18],layer1[20],amt[1]);
mux_2x1 L2_19(layer2[19],layer1[19],layer1[21],amt[1]);
mux_2x1 L2_20(layer2[20],layer1[20],layer1[22],amt[1]);
mux_2x1 L2_21(layer2[21],layer1[21],layer1[23],amt[1]);
mux_2x1 L2_22(layer2[22],layer1[22],layer1[24],amt[1]);
mux_2x1 L2_23(layer2[23],layer1[23],layer1[25],amt[1]);
mux_2x1 L2_24(layer2[24],layer1[24],layer1[26],amt[1]);
mux_2x1 L2_25(layer2[25],layer1[25],layer1[27],amt[1]);
mux_2x1 L2_26(layer2[26],layer1[26],layer1[28],amt[1]);
mux_2x1 L2_27(layer2[27],layer1[27],layer1[29],amt[1]);
mux_2x1 L2_28(layer2[28],layer1[28],layer1[30],amt[1]);
mux_2x1 L2_29(layer2[29],layer1[29],layer1[31],amt[1]);
mux_2x1 L2_30(layer2[30],layer1[30],empty,amt[1]);
mux_2x1 L2_31(layer2[31],layer1[31],empty,amt[1]);
mux_2x1 L3_0(layer3[0],layer2[0],layer2[4],amt[2]);
mux_2x1 L3_1(layer3[1],layer2[1],layer2[5],amt[2]);
mux_2x1 L3_2(layer3[2],layer2[2],layer2[6],amt[2]);
mux_2x1 L3_3(layer3[3],layer2[3],layer2[7],amt[2]);
mux_2x1 L3_4(layer3[4],layer2[4],layer2[8],amt[2]);
mux_2x1 L3_5(layer3[5],layer2[5],layer2[9],amt[2]);
mux_2x1 L3_6(layer3[6],layer2[6],layer2[10],amt[2]);
mux_2x1 L3_7(layer3[7],layer2[7],layer2[11],amt[2]);
mux_2x1 L3_8(layer3[8],layer2[8],layer2[12],amt[2]);
mux_2x1 L3_9(layer3[9],layer2[9],layer2[13],amt[2]);
mux_2x1 L3_10(layer3[10],layer2[10],layer2[14],amt[2]);
mux_2x1 L3_11(layer3[11],layer2[11],layer2[15],amt[2]);
mux_2x1 L3_12(layer3[12],layer2[12],layer2[16],amt[2]);
mux_2x1 L3_13(layer3[13],layer2[13],layer2[17],amt[2]);
mux_2x1 L3_14(layer3[14],layer2[14],layer2[18],amt[2]);
mux_2x1 L3_15(layer3[15],layer2[15],layer2[19],amt[2]);
mux_2x1 L3_16(layer3[16],layer2[16],layer2[20],amt[2]);
mux_2x1 L3_17(layer3[17],layer2[17],layer2[21],amt[2]);
mux_2x1 L3_18(layer3[18],layer2[18],layer2[22],amt[2]);
mux_2x1 L3_19(layer3[19],layer2[19],layer2[23],amt[2]);
mux_2x1 L3_20(layer3[20],layer2[20],layer2[24],amt[2]);
mux_2x1 L3_21(layer3[21],layer2[21],layer2[25],amt[2]);
mux_2x1 L3_22(layer3[22],layer2[22],layer2[26],amt[2]);
mux_2x1 L3_23(layer3[23],layer2[23],layer2[27],amt[2]);
mux_2x1 L3_24(layer3[24],layer2[24],layer2[28],amt[2]);
mux_2x1 L3_25(layer3[25],layer2[25],layer2[29],amt[2]);
mux_2x1 L3_26(layer3[26],layer2[26],layer2[30],amt[2]);
mux_2x1 L3_27(layer3[27],layer2[27],layer2[31],amt[2]);
mux_2x1 L3_28(layer3[28],layer2[28],empty,amt[2]);
mux_2x1 L3_29(layer3[29],layer2[29],empty,amt[2]);
mux_2x1 L3_30(layer3[30],layer2[30],empty,amt[2]);
mux_2x1 L3_31(layer3[31],layer2[31],empty,amt[2]);
mux_2x1 L4_0(layer4[0],layer3[0],layer3[8],amt[3]);
mux_2x1 L4_1(layer4[1],layer3[1],layer3[9],amt[3]);
mux_2x1 L4_2(layer4[2],layer3[2],layer3[10],amt[3]);
mux_2x1 L4_3(layer4[3],layer3[3],layer3[11],amt[3]);
mux_2x1 L4_4(layer4[4],layer3[4],layer3[12],amt[3]);
mux_2x1 L4_5(layer4[5],layer3[5],layer3[13],amt[3]);
mux_2x1 L4_6(layer4[6],layer3[6],layer3[14],amt[3]);
mux_2x1 L4_7(layer4[7],layer3[7],layer3[15],amt[3]);
mux_2x1 L4_8(layer4[8],layer3[8],layer3[16],amt[3]);
mux_2x1 L4_9(layer4[9],layer3[9],layer3[17],amt[3]);
mux_2x1 L4_10(layer4[10],layer3[10],layer3[18],amt[3]);
mux_2x1 L4_11(layer4[11],layer3[11],layer3[19],amt[3]);
mux_2x1 L4_12(layer4[12],layer3[12],layer3[20],amt[3]);
mux_2x1 L4_13(layer4[13],layer3[13],layer3[21],amt[3]);
mux_2x1 L4_14(layer4[14],layer3[14],layer3[22],amt[3]);
mux_2x1 L4_15(layer4[15],layer3[15],layer3[23],amt[3]);
mux_2x1 L4_16(layer4[16],layer3[16],layer3[24],amt[3]);
mux_2x1 L4_17(layer4[17],layer3[17],layer3[25],amt[3]);
mux_2x1 L4_18(layer4[18],layer3[18],layer3[26],amt[3]);
mux_2x1 L4_19(layer4[19],layer3[19],layer3[27],amt[3]);
mux_2x1 L4_20(layer4[20],layer3[20],layer3[28],amt[3]);
mux_2x1 L4_21(layer4[21],layer3[21],layer3[29],amt[3]);
mux_2x1 L4_22(layer4[22],layer3[22],layer3[30],amt[3]);
mux_2x1 L4_23(layer4[23],layer3[23],layer3[31],amt[3]);
mux_2x1 L4_24(layer4[24],layer3[24],empty,amt[3]);
mux_2x1 L4_25(layer4[25],layer3[25],empty,amt[3]);
mux_2x1 L4_26(layer4[26],layer3[26],empty,amt[3]);
mux_2x1 L4_27(layer4[27],layer3[27],empty,amt[3]);
mux_2x1 L4_28(layer4[28],layer3[28],empty,amt[3]);
mux_2x1 L4_29(layer4[29],layer3[29],empty,amt[3]);
mux_2x1 L4_30(layer4[30],layer3[30],empty,amt[3]);
mux_2x1 L4_31(layer4[31],layer3[31],empty,amt[3]);
mux_2x1 L5_0(layer5[0],layer4[0],layer4[16],amt[4]);
mux_2x1 L5_1(layer5[1],layer4[1],layer4[17],amt[4]);
mux_2x1 L5_2(layer5[2],layer4[2],layer4[18],amt[4]);
mux_2x1 L5_3(layer5[3],layer4[3],layer4[19],amt[4]);
mux_2x1 L5_4(layer5[4],layer4[4],layer4[20],amt[4]);
mux_2x1 L5_5(layer5[5],layer4[5],layer4[21],amt[4]);
mux_2x1 L5_6(layer5[6],layer4[6],layer4[22],amt[4]);
mux_2x1 L5_7(layer5[7],layer4[7],layer4[23],amt[4]);
mux_2x1 L5_8(layer5[8],layer4[8],layer4[24],amt[4]);
mux_2x1 L5_9(layer5[9],layer4[9],layer4[25],amt[4]);
mux_2x1 L5_10(layer5[10],layer4[10],layer4[26],amt[4]);
mux_2x1 L5_11(layer5[11],layer4[11],layer4[27],amt[4]);
mux_2x1 L5_12(layer5[12],layer4[12],layer4[28],amt[4]);
mux_2x1 L5_13(layer5[13],layer4[13],layer4[29],amt[4]);
mux_2x1 L5_14(layer5[14],layer4[14],layer4[30],amt[4]);
mux_2x1 L5_15(layer5[15],layer4[15],layer4[31],amt[4]);
mux_2x1 L5_16(layer5[16],layer4[16],empty,amt[4]);
mux_2x1 L5_17(layer5[17],layer4[17],empty,amt[4]);
mux_2x1 L5_18(layer5[18],layer4[18],empty,amt[4]);
mux_2x1 L5_19(layer5[19],layer4[19],empty,amt[4]);
mux_2x1 L5_20(layer5[20],layer4[20],empty,amt[4]);
mux_2x1 L5_21(layer5[21],layer4[21],empty,amt[4]);
mux_2x1 L5_22(layer5[22],layer4[22],empty,amt[4]);
mux_2x1 L5_23(layer5[23],layer4[23],empty,amt[4]);
mux_2x1 L5_24(layer5[24],layer4[24],empty,amt[4]);
mux_2x1 L5_25(layer5[25],layer4[25],empty,amt[4]);
mux_2x1 L5_26(layer5[26],layer4[26],empty,amt[4]);
mux_2x1 L5_27(layer5[27],layer4[27],empty,amt[4]);
mux_2x1 L5_28(layer5[28],layer4[28],empty,amt[4]);
mux_2x1 L5_29(layer5[29],layer4[29],empty,amt[4]);
mux_2x1 L5_30(layer5[30],layer4[30],empty,amt[4]);
mux_2x1 L5_31(layer5[31],layer4[31],empty,amt[4]);

mux_2x1 F0(out[0],layer5[0],layer5[31],rev);
mux_2x1 F1(out[1],layer5[1],layer5[30],rev);
mux_2x1 F2(out[2],layer5[2],layer5[29],rev);
mux_2x1 F3(out[3],layer5[3],layer5[28],rev);
mux_2x1 F4(out[4],layer5[4],layer5[27],rev);
mux_2x1 F5(out[5],layer5[5],layer5[26],rev);
mux_2x1 F6(out[6],layer5[6],layer5[25],rev);
mux_2x1 F7(out[7],layer5[7],layer5[24],rev);
mux_2x1 F8(out[8],layer5[8],layer5[23],rev);
mux_2x1 F9(out[9],layer5[9],layer5[22],rev);
mux_2x1 F10(out[10],layer5[10],layer5[21],rev);
mux_2x1 F11(out[11],layer5[11],layer5[20],rev);
mux_2x1 F12(out[12],layer5[12],layer5[19],rev);
mux_2x1 F13(out[13],layer5[13],layer5[18],rev);
mux_2x1 F14(out[14],layer5[14],layer5[17],rev);
mux_2x1 F15(out[15],layer5[15],layer5[16],rev);
mux_2x1 F16(out[16],layer5[16],layer5[15],rev);
mux_2x1 F17(out[17],layer5[17],layer5[14],rev);
mux_2x1 F18(out[18],layer5[18],layer5[13],rev);
mux_2x1 F19(out[19],layer5[19],layer5[12],rev);
mux_2x1 F20(out[20],layer5[20],layer5[11],rev);
mux_2x1 F21(out[21],layer5[21],layer5[10],rev);
mux_2x1 F22(out[22],layer5[22],layer5[9],rev);
mux_2x1 F23(out[23],layer5[23],layer5[8],rev);
mux_2x1 F24(out[24],layer5[24],layer5[7],rev);
mux_2x1 F25(out[25],layer5[25],layer5[6],rev);
mux_2x1 F26(out[26],layer5[26],layer5[5],rev);
mux_2x1 F27(out[27],layer5[27],layer5[4],rev);
mux_2x1 F28(out[28],layer5[28],layer5[3],rev);
mux_2x1 F29(out[29],layer5[29],layer5[2],rev);
mux_2x1 F30(out[30],layer5[30],layer5[1],rev);
mux_2x1 F31(out[31],layer5[31],layer5[0],rev);
endmodule