module extend(output[31:0] zero,output[31:0] sign,input[15:0] imm);

buf b31  (zero[31],1'b0);
buf b30  (zero[30],1'b0);
buf b29  (zero[29],1'b0);
buf b28  (zero[28],1'b0);
buf b27  (zero[27],1'b0);
buf b26  (zero[26],1'b0);
buf b25  (zero[25],1'b0);
buf b24  (zero[24],1'b0);
buf b23  (zero[23],1'b0);
buf b22  (zero[22],1'b0);
buf b21  (zero[21],1'b0);
buf b20  (zero[20],1'b0);
buf b19  (zero[19],1'b0);
buf b18  (zero[18],1'b0);
buf b17  (zero[17],1'b0);
buf b16  (zero[16],1'b0);
buf b15  (zero[15],imm[15]);
buf b14  (zero[14],imm[14]);
buf b13  (zero[13],imm[13]);
buf b12  (zero[12],imm[12]);
buf b11  (zero[11],imm[11]);
buf b10  (zero[10],imm[10]);
buf b9  (zero[9],imm[9]);
buf b8  (zero[8],imm[8]);
buf b7  (zero[7],imm[7]);
buf b6  (zero[6],imm[6]);
buf b5  (zero[5],imm[5]);
buf b4  (zero[4],imm[4]);
buf b3  (zero[3],imm[3]);
buf b2  (zero[2],imm[2]);
buf b1  (zero[1],imm[1]);
buf b0  (zero[0],imm[0]);

buf bb31  (sign[31],imm[15]);
buf bb30  (sign[30],imm[15]);
buf bb29  (sign[29],imm[15]);
buf bb28  (sign[28],imm[15]);
buf bb27  (sign[27],imm[15]);
buf bb26  (sign[26],imm[15]);
buf bb25  (sign[25],imm[15]);
buf bb24  (sign[24],imm[15]);
buf bb23  (sign[23],imm[15]);
buf bb22  (sign[22],imm[15]);
buf bb21  (sign[21],imm[15]);
buf bb20  (sign[20],imm[15]);
buf bb19  (sign[19],imm[15]);
buf bb18  (sign[18],imm[15]);
buf bb17  (sign[17],imm[15]);
buf bb16  (sign[16],imm[15]);
buf bb15  (sign[15],imm[15]);
buf bb14  (sign[14],imm[14]);
buf bb13  (sign[13],imm[13]);
buf bb12  (sign[12],imm[12]);
buf bb11  (sign[11],imm[11]);
buf bb10  (sign[10],imm[10]);
buf bb9  (sign[9],imm[9]);
buf bb8  (sign[8],imm[8]);
buf bb7  (sign[7],imm[7]);
buf bb6  (sign[6],imm[6]);
buf bb5  (sign[5],imm[5]);
buf bb4  (sign[4],imm[4]);
buf bb3  (sign[3],imm[3]);
buf bb2  (sign[2],imm[2]);
buf bb1  (sign[1],imm[1]);
buf bb0  (sign[0],imm[0]);


endmodule